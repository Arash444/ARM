module ARM (clk, rst);
    
    input clk, rst;

endmodule