module Cache_cntrlr (
    
);
    
endmodule