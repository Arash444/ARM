module Instru_mem (
    addr,
    instru
);

    input [31:0] addr;
    output reg [31:0] instru;

    always @(addr) begin
        case(addr)
            32'd0: instru = 32'b1110_00_1_1101_0_0000_0000_000000010100;
            32'd4: instru = 32'b1110_00_1_1101_0_0000_0001_101000000001;            
            32'd8: instru = 32'b1110_00_1_1101_0_0000_0010_000100000011;           
            32'd12: instru = 32'b1110_00_0_0100_1_0010_0011_000000000010;            
            32'd16: instru = 32'b1110_00_0_0101_0_0000_0100_000000000000;            
            32'd20: instru = 32'b1110_00_0_0010_0_0100_0101_000100000100;           
            32'd24: instru = 32'b1110_00_0_0110_0_0000_0110_000010100000;           
            32'd28: instru = 32'b1110_00_0_1100_0_0101_0111_000101000010;            
            32'd32: instru = 32'b1110_00_0_0000_0_0111_1000_000000000011;           
            32'd36: instru = 32'b1110_00_0_1111_0_0000_1001_000000000110;
            32'd40: instru = 32'b1110_00_0_0001_0_0100_1010_000000000101;
            32'd44: instru = 32'b1110_00_0_1010_1_1000_0000_000000000110; 
            32'd48: instru = 32'b0001_00_0_0100_0_0001_0001_000000000001;
            32'd52: instru = 32'b1110_00_0_1000_1_1001_0000_000000001000;
            32'd56: instru = 32'b0000_00_0_0100_0_0010_0010_000000000010;
            32'd60: instru = 32'b1110_00_1_1101_0_0000_0000_101100000001;
            32'd64: instru = 32'b1110_01_0_0100_0_0000_0001_000000000000;
            32'd68: instru = 32'b1110_01_0_0100_1_0000_1011_000000000000;
            32'd72: instru = 32'b1110_01_0_0100_0_0000_0010_000000000100;
            32'd76: instru = 32'b1110_01_0_0100_0_0000_0011_000000001000; 
            32'd80: instru = 32'b1110_01_0_0100_0_0000_0100_000000001101; 
            32'd84: instru = 32'b1110_01_0_0100_0_0000_0101_000000010000; 
            32'd88: instru = 32'b1110_01_0_0100_0_0000_0110_000000010100; 
            32'd92: instru = 32'b1110_01_0_0100_1_0000_1010_000000000100; 
            32'd96: instru = 32'b1110_01_0_0100_0_0000_0111_000000011000; 
            32'd100: instru = 32'b1110_00_1_1101_0_0000_0001_000000000100; 
            32'd104: instru = 32'b1110_00_1_1101_0_0000_0010_000000000000; 
            32'd108: instru = 32'b1110_00_1_1101_0_0000_0011_000000000000; 
            32'd112: instru = 32'b1110_00_0_0100_0_0000_0100_000100000011; 	
            32'd116: instru = 32'b1110_01_0_0100_1_0100_0101_000000000000; 
            32'd120: instru = 32'b1110_01_0_0100_1_0100_0110_000000000100; 
            32'd124: instru = 32'b1110_00_0_1010_1_0101_0000_000000000110; 
            32'd128: instru = 32'b1100_01_0_0100_0_0100_0110_000000000000; 
            32'd132: instru = 32'b1100_01_0_0100_0_0100_0101_000000000100; 
            32'd136: instru = 32'b1110_00_1_0100_0_0011_0011_000000000001; 
            32'd140: instru = 32'b1110_00_1_1010_1_0011_0000_000000000011; 
            32'd144: instru = 32'b1011_10_1_0_111111111111111111110111; 
            32'd148: instru = 32'b1110_00_1_0100_0_0010_0010_000000000001; 
            32'd152: instru = 32'b1110_00_0_1010_1_0010_0000_000000000001; 
            32'd156: instru = 32'b1011_10_1_0_111111111111111111110011; 
            32'd160: instru = 32'b1110_01_0_0100_1_0000_0001_000000000000; 
            32'd164: instru = 32'b1110_01_0_0100_1_0000_0010_000000000100; 
            32'd168: instru = 32'b1110_01_0_0100_1_0000_0011_000000001000; 
            32'd172: instru = 32'b1110_01_0_0100_1_0000_0100_000000001100; 
            32'd176: instru = 32'b1110_01_0_0100_1_0000_0101_000000010000; 
            32'd180: instru = 32'b1110_01_0_0100_1_0000_0110_000000010100; 
            32'd184: instru = 32'b1110_10_1_0_111111111111111111111111;
            default: instru = 32'b0;
        endcase
    end

endmodule